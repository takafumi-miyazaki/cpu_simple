module instruction_memory(A, B);
   input [3:0] A;
   output [7:0] B;
   reg [7:0] 	im[15:0];

   
   
endmodule // instruction_memory
